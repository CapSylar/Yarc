package riscv_pkg;



endpackage: riscv_pkg